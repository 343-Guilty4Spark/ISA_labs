package constants is
    constant Nbit : integer := 7;
end package;